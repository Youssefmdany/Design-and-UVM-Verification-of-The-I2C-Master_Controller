


package I2C_pkg;


 import uvm_pkg::*;
 
 `include "uvm_macros.svh"
  
  
  `include "I2C_seq_item.sv"
  `include "Sequence.sv"
  `include "Sequencer.sv"   
  `include "Driver.sv"  
  `include "Monitor.sv"
  `include "Agent.sv"  
  `include "Scoreboard.sv"
  `include "Environment.sv"  
  `include "I2C_Test.sv"

 

endpackage 